`define ALU_TYPE 8
`define ALU_ADD 0
`define ALU_SLT 1
`define ALU_SLL 2
`define ALU_SRL 3
`define ALU_SRA 4
`define ALU_XOR 5
`define ALU_OR  6
`define ALU_AND 7

