module ps2_top_apb(
  input         clock,
  input         reset,
  input  [31:0] in_paddr,
  input         in_psel,
  input         in_penable,
  input  [2:0]  in_pprot,
  input         in_pwrite,
  input  [31:0] in_pwdata,
  input  [3:0]  in_pstrb,
  output        in_pready,
  output [31:0] in_prdata,
  output        in_pslverr,

  input         ps2_clk,
  input         ps2_data
);

reg in_ready, ready;

assign in_pready = in_ready;
always@(posedge clock)begin
  if(in_penable && !in_ready)
    in_ready <= 1;
  else if(in_ready)
    in_ready <= 0;
  end

reg [9:0] buffer;        // ps2_data bits
reg [7:0] fifo[7:0];     // data fifo
reg [2:0] w_ptr,r_ptr;   // fifo write and read pointers
reg [3:0] count;  // count ps2_data bits
// detect falling edge of ps2_clk
reg [2:0] ps2_clk_sync;

always @(posedge clock) begin
  ps2_clk_sync <=  {ps2_clk_sync[1:0],ps2_clk};
end

wire sampling = ps2_clk_sync[2] & ~ps2_clk_sync[1];

always @(posedge clock) begin
  if (reset) begin // reset
    count <= 0; w_ptr <= 0; r_ptr <= 0; ready<= 0;
  end
  else begin
    if ( ready ) begin // read to output next data
      if(in_ready) //read next data
      begin
          r_ptr <= r_ptr + 3'b1;
          fifo[r_ptr] <= 0;
          if(w_ptr==(r_ptr+1'b1)) //empty
              ready <= 1'b0;
      end
    end
    if (sampling) begin
      if (count == 4'd10) begin
        if ((buffer[0] == 0) &&  // start bit
          (ps2_data)       &&  // stop bit
          (^buffer[9:1])) begin      // odd  parity
          fifo[w_ptr] <= buffer[8:1];  // kbd scan code
          w_ptr <= w_ptr+3'b1;
          ready <= 1'b1;
          //$display("receive %x", buffer[8:1]);
        end
        count <= 0;     // for next
      end else begin
        buffer[count] <= ps2_data;  // store ps2_data
        count <= count + 3'b1;
      end
    end
  end
end
assign in_prdata = {24'b0, fifo[r_ptr]};


endmodule
