
`define BRANCH_MID 7:0
`define BRANCH 0
`define BRANCH_BACK 1
`define BEQ 2
`define ZERO 3
`define BNE 4
`define BLT 5
`define CMP 6
`define BGE 7

